module drive_one( output one );

// Insert your code here
    assign one = 1'b1;

endmodule